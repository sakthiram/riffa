library verilog;
use verilog.vl_types.all;
entity channel_128 is
    generic(
        C_DATA_WIDTH    : vl_logic_vector(0 to 8) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        C_MAX_READ_REQ  : integer := 2;
        C_RX_FIFO_DEPTH : integer := 1024;
        C_TX_FIFO_DEPTH : integer := 512;
        C_SG_FIFO_DEPTH : integer := 1024;
        C_DATA_WORD_WIDTH: vl_notype
    );
    port(
        CLK             : in     vl_logic;
        RST             : in     vl_logic;
        CONFIG_MAX_READ_REQUEST_SIZE: in     vl_logic_vector(2 downto 0);
        CONFIG_MAX_PAYLOAD_SIZE: in     vl_logic_vector(2 downto 0);
        PIO_DATA        : in     vl_logic_vector(31 downto 0);
        ENG_DATA        : in     vl_logic_vector;
        SG_RX_BUF_RECVD : out    vl_logic;
        SG_RX_BUF_LEN_VALID: in     vl_logic;
        SG_RX_BUF_ADDR_HI_VALID: in     vl_logic;
        SG_RX_BUF_ADDR_LO_VALID: in     vl_logic;
        SG_TX_BUF_RECVD : out    vl_logic;
        SG_TX_BUF_LEN_VALID: in     vl_logic;
        SG_TX_BUF_ADDR_HI_VALID: in     vl_logic;
        SG_TX_BUF_ADDR_LO_VALID: in     vl_logic;
        TXN_RX_LEN_VALID: in     vl_logic;
        TXN_RX_OFF_LAST_VALID: in     vl_logic;
        TXN_RX_DONE_LEN : out    vl_logic_vector(31 downto 0);
        TXN_RX_DONE     : out    vl_logic;
        TXN_RX_DONE_ACK : in     vl_logic;
        TXN_TX          : out    vl_logic;
        TXN_TX_ACK      : in     vl_logic;
        TXN_TX_LEN      : out    vl_logic_vector(31 downto 0);
        TXN_TX_OFF_LAST : out    vl_logic_vector(31 downto 0);
        TXN_TX_DONE_LEN : out    vl_logic_vector(31 downto 0);
        TXN_TX_DONE     : out    vl_logic;
        TXN_TX_DONE_ACK : in     vl_logic;
        RX_REQ          : out    vl_logic;
        RX_REQ_ACK      : in     vl_logic;
        RX_REQ_TAG      : out    vl_logic_vector(1 downto 0);
        RX_REQ_ADDR     : out    vl_logic_vector(63 downto 0);
        RX_REQ_LEN      : out    vl_logic_vector(9 downto 0);
        TX_REQ          : out    vl_logic;
        TX_REQ_ACK      : in     vl_logic;
        TX_ADDR         : out    vl_logic_vector(63 downto 0);
        TX_LEN          : out    vl_logic_vector(9 downto 0);
        TX_DATA         : out    vl_logic_vector;
        TX_DATA_REN     : in     vl_logic;
        TX_SENT         : in     vl_logic;
        MAIN_DATA_EN    : in     vl_logic_vector;
        MAIN_DONE       : in     vl_logic;
        MAIN_ERR        : in     vl_logic;
        SG_RX_DATA_EN   : in     vl_logic_vector;
        SG_RX_DONE      : in     vl_logic;
        SG_RX_ERR       : in     vl_logic;
        SG_TX_DATA_EN   : in     vl_logic_vector;
        SG_TX_DONE      : in     vl_logic;
        SG_TX_ERR       : in     vl_logic;
        CHNL_RX_CLK     : in     vl_logic;
        CHNL_RX         : out    vl_logic;
        CHNL_RX_ACK     : in     vl_logic;
        CHNL_RX_LAST    : out    vl_logic;
        CHNL_RX_LEN     : out    vl_logic_vector(31 downto 0);
        CHNL_RX_OFF     : out    vl_logic_vector(30 downto 0);
        CHNL_RX_DATA    : out    vl_logic_vector;
        CHNL_RX_DATA_VALID: out    vl_logic;
        CHNL_RX_DATA_REN: in     vl_logic;
        CHNL_TX_CLK     : in     vl_logic;
        CHNL_TX         : in     vl_logic;
        CHNL_TX_ACK     : out    vl_logic;
        CHNL_TX_LAST    : in     vl_logic;
        CHNL_TX_LEN     : in     vl_logic_vector(31 downto 0);
        CHNL_TX_OFF     : in     vl_logic_vector(30 downto 0);
        CHNL_TX_DATA    : in     vl_logic_vector;
        CHNL_TX_DATA_VALID: in     vl_logic;
        CHNL_TX_DATA_REN: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_MAX_READ_REQ : constant is 1;
    attribute mti_svvh_generic_type of C_RX_FIFO_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of C_TX_FIFO_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of C_SG_FIFO_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of C_DATA_WORD_WIDTH : constant is 3;
end channel_128;
