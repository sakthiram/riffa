`include "functions.vh"
`define DATA_WIDTH 10'd256
`define DATA_WORD_WIDTH clog2((`DATA_WIDTH/32)+1)
